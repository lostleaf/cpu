module test;
always begin
	#10
	#10 $finish;
end
endmodule