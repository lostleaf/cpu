module data_memory_testbench ;
    `include "parameters.v"
endmodule