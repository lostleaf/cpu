module def_param;
	defparam 
	CPU.alu_rs[0].fuindex = 0,
	CPU.alu_rs[1].fuindex = 1,
	CPU.alu_rs[2].fuindex = 2;
endmodule