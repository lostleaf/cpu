module rs ();
    
endmodule