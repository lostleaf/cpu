module inst_decode (inst, reg1, reg2, out_alu1, out_alu2, decode_enable);
    input wire [WORD_SIZE-1:0] inst, reg1, reg2;

endmodule